----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:34:35 08/22/2019 
-- Design Name: 
-- Module Name:    myFFDR - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity myFFDR is
port(clk: in std_logic;
		rst: in std_logic;
		d: in std_logic;
		q: out std_logic);
end myFFDR;

architecture Arch_myFFDR of myFFDR is

begin

process(clk)
begin
	if(rising_edge(clk)) then
		if(rst = '1') then
				q <= '0';
			else
				q <= d;
		end if;
	end if;
end process;
	
end Arch_myFFDR;

